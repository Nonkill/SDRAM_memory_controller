module memory_controller(
    port_list
);
    
endmodule